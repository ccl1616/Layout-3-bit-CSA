* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT MA_MOS
** N=9 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV gnd inv_in vdd inv_out
** N=4 EP=4 IP=0 FDC=2
M0 inv_out inv_in gnd gnd N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06 $X=1260 $Y=220 $D=0
M1 inv_out inv_in vdd vdd P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06 $X=1260 $Y=1660 $D=1
.ENDS
***************************************
.SUBCKT FA GND VDD a b c_in sum c_out
** N=20 EP=7 IP=24 FDC=28
M0 10 a GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=1170 $Y=1510 $D=0
M1 GND b 10 GND N_18 L=1.8e-07 W=4.7e-07 AD=3.055e-13 AS=1.6685e-13 PD=1.3e-06 PS=7.1e-07 $X=1170 $Y=2400 $D=0
M2 10 c_in GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.7155e-13 AS=3.055e-13 PD=7.3e-07 PS=1.3e-06 $X=1170 $Y=3290 $D=0
M3 8 9 10 GND N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.7155e-13 PD=1.45e-06 PS=7.3e-07 $X=1170 $Y=4200 $D=0
M4 18 a GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=1940 $Y=1510 $D=0
M5 19 b 18 GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=1.6685e-13 PD=7.1e-07 PS=7.1e-07 $X=1940 $Y=2400 $D=0
M6 8 c_in 19 GND N_18 L=1.8e-07 W=4.7e-07 AD=2.867e-13 AS=1.6685e-13 PD=1.69e-06 PS=7.1e-07 $X=1940 $Y=3290 $D=0
M7 20 a GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=2730 $Y=1510 $D=0
M8 9 b 20 GND N_18 L=1.8e-07 W=4.7e-07 AD=2.773e-13 AS=1.6685e-13 PD=1.65e-06 PS=7.1e-07 $X=2730 $Y=2400 $D=0
M9 GND a 11 GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=3510 $Y=1510 $D=0
M10 11 b GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=1.6685e-13 PD=7.1e-07 PS=7.1e-07 $X=3510 $Y=2400 $D=0
M11 9 c_in 11 GND N_18 L=1.8e-07 W=4.7e-07 AD=2.867e-13 AS=1.6685e-13 PD=1.69e-06 PS=7.1e-07 $X=3510 $Y=3290 $D=0
M12 VDD a 13 VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=5140 $Y=1510 $D=1
M13 13 b VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=1.6685e-13 PD=7.1e-07 PS=7.1e-07 $X=5140 $Y=2400 $D=1
M14 9 c_in 13 VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.867e-13 AS=1.6685e-13 PD=1.69e-06 PS=7.1e-07 $X=5140 $Y=3290 $D=1
M15 15 a VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=5920 $Y=1510 $D=1
M16 9 b 15 VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.773e-13 AS=1.6685e-13 PD=1.65e-06 PS=7.1e-07 $X=5920 $Y=2400 $D=1
M17 16 a VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=6710 $Y=1510 $D=1
M18 17 b 16 VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=1.6685e-13 PD=7.1e-07 PS=7.1e-07 $X=6710 $Y=2400 $D=1
M19 8 c_in 17 VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.867e-13 AS=1.6685e-13 PD=1.69e-06 PS=7.1e-07 $X=6710 $Y=3290 $D=1
M20 12 a VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=7480 $Y=1510 $D=1
M21 VDD b 12 VDD P_18 L=1.8e-07 W=4.7e-07 AD=3.055e-13 AS=1.6685e-13 PD=1.3e-06 PS=7.1e-07 $X=7480 $Y=2400 $D=1
M22 12 c_in VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.7155e-13 AS=3.055e-13 PD=7.3e-07 PS=1.3e-06 $X=7480 $Y=3290 $D=1
M23 8 9 12 VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.7155e-13 PD=1.45e-06 PS=7.3e-07 $X=7480 $Y=4200 $D=1
X26 GND 8 VDD sum INV $T=11740 3620 1 270 $X=9110 $Y=1190
X27 GND 9 VDD c_out INV $T=11740 2940 0 90 $X=9110 $Y=3210
.ENDS
***************************************
.SUBCKT MUX21 ctrl GND VDD in2 out in1
** N=7 EP=6 IP=0 FDC=6
M0 7 ctrl GND GND N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=2.303e-13 PD=1.49e-06 PS=1.45e-06 $X=2190 $Y=380 $D=0
M1 out ctrl in2 GND N_18 L=1.8e-07 W=4.7e-07 AD=1.222e-13 AS=2.35e-13 PD=5.2e-07 PS=1.47e-06 $X=3800 $Y=380 $D=0
M2 in1 7 out GND N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.222e-13 PD=1.45e-06 PS=5.2e-07 $X=4500 $Y=380 $D=0
M3 7 ctrl VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=2.303e-13 PD=1.49e-06 PS=1.45e-06 $X=2190 $Y=2460 $D=1
M4 out 7 in2 VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.222e-13 AS=2.35e-13 PD=5.2e-07 PS=1.47e-06 $X=3800 $Y=2460 $D=1
M5 in1 ctrl out VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.222e-13 PD=1.45e-06 PS=5.2e-07 $X=4500 $Y=2460 $D=1
.ENDS
***************************************
.SUBCKT ADDER3 B0 GND A0 A1 B1 VDD A2 B2 CIN S0 S1 S2 COUT
** N=25 EP=13 IP=66 FDC=192
X0 GND VDD A0 B0 GND 20 9 FA $T=-10 0 0 0 $X=0 $Y=0
X1 GND VDD A1 B1 9 21 10 FA $T=-10 5410 0 0 $X=0 $Y=5410
X2 GND VDD A2 B2 10 22 11 FA $T=-10 10820 0 0 $X=0 $Y=10820
X3 GND VDD A0 B0 VDD 23 13 FA $T=28460 10 1 180 $X=16240 $Y=10
X4 GND VDD A1 B1 13 24 14 FA $T=28460 5420 1 180 $X=16240 $Y=5420
X5 GND VDD A2 B2 14 25 12 FA $T=28460 10830 1 180 $X=16240 $Y=10830
X6 CIN GND VDD 23 S0 20 MUX21 $T=12190 6790 0 270 $X=12190 $Y=970
X7 CIN GND VDD 24 S1 21 MUX21 $T=12190 12020 0 270 $X=12190 $Y=6200
X8 CIN GND VDD 25 S2 22 MUX21 $T=12190 17250 0 270 $X=12190 $Y=11430
X9 CIN GND VDD 12 COUT 11 MUX21 $T=12190 22480 0 270 $X=12190 $Y=16660
.ENDS
***************************************
