* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT MA_MOS
** N=9 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV gnd inv_in vdd inv_out
** N=4 EP=4 IP=0 FDC=2
M0 inv_out inv_in gnd gnd N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06 $X=1260 $Y=220 $D=0
M1 inv_out inv_in vdd vdd P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06 $X=1260 $Y=1660 $D=1
.ENDS
***************************************
.SUBCKT FA GND VDD a b c_in sum c_out
** N=20 EP=7 IP=24 FDC=28
M0 9 a GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=1870 $Y=1510 $D=0
M1 GND b 9 GND N_18 L=1.8e-07 W=4.7e-07 AD=3.055e-13 AS=1.6685e-13 PD=1.3e-06 PS=7.1e-07 $X=1870 $Y=2400 $D=0
M2 9 c_in GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.7155e-13 AS=3.055e-13 PD=7.3e-07 PS=1.3e-06 $X=1870 $Y=3290 $D=0
M3 3 7 9 GND N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.7155e-13 PD=1.45e-06 PS=7.3e-07 $X=1870 $Y=4200 $D=0
M4 18 a GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=2640 $Y=1510 $D=0
M5 19 b 18 GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=1.6685e-13 PD=7.1e-07 PS=7.1e-07 $X=2640 $Y=2400 $D=0
M6 3 c_in 19 GND N_18 L=1.8e-07 W=4.7e-07 AD=2.867e-13 AS=1.6685e-13 PD=1.69e-06 PS=7.1e-07 $X=2640 $Y=3290 $D=0
M7 20 a GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=3430 $Y=1510 $D=0
M8 7 b 20 GND N_18 L=1.8e-07 W=4.7e-07 AD=2.773e-13 AS=1.6685e-13 PD=1.65e-06 PS=7.1e-07 $X=3430 $Y=2400 $D=0
M9 GND a 10 GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=4210 $Y=1510 $D=0
M10 10 b GND GND N_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=1.6685e-13 PD=7.1e-07 PS=7.1e-07 $X=4210 $Y=2400 $D=0
M11 7 c_in 10 GND N_18 L=1.8e-07 W=4.7e-07 AD=2.867e-13 AS=1.6685e-13 PD=1.69e-06 PS=7.1e-07 $X=4210 $Y=3290 $D=0
M12 VDD a 12 VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=5840 $Y=1510 $D=1
M13 12 b VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=1.6685e-13 PD=7.1e-07 PS=7.1e-07 $X=5840 $Y=2400 $D=1
M14 7 c_in 12 VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.867e-13 AS=1.6685e-13 PD=1.69e-06 PS=7.1e-07 $X=5840 $Y=3290 $D=1
M15 15 a VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=6620 $Y=1510 $D=1
M16 7 b 15 VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.773e-13 AS=1.6685e-13 PD=1.65e-06 PS=7.1e-07 $X=6620 $Y=2400 $D=1
M17 16 a VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=7410 $Y=1510 $D=1
M18 17 b 16 VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=1.6685e-13 PD=7.1e-07 PS=7.1e-07 $X=7410 $Y=2400 $D=1
M19 3 c_in 17 VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.867e-13 AS=1.6685e-13 PD=1.69e-06 PS=7.1e-07 $X=7410 $Y=3290 $D=1
M20 11 a VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.6685e-13 AS=2.303e-13 PD=7.1e-07 PS=1.45e-06 $X=8180 $Y=1510 $D=1
M21 VDD b 11 VDD P_18 L=1.8e-07 W=4.7e-07 AD=3.055e-13 AS=1.6685e-13 PD=1.3e-06 PS=7.1e-07 $X=8180 $Y=2400 $D=1
M22 11 c_in VDD VDD P_18 L=1.8e-07 W=4.7e-07 AD=1.7155e-13 AS=3.055e-13 PD=7.3e-07 PS=1.3e-06 $X=8180 $Y=3290 $D=1
M23 3 7 11 VDD P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.7155e-13 PD=1.45e-06 PS=7.3e-07 $X=8180 $Y=4200 $D=1
X26 GND 3 VDD sum INV $T=12440 3620 1 270 $X=9810 $Y=1190
X27 GND 7 VDD c_out INV $T=12440 2940 0 90 $X=9810 $Y=3210
.ENDS
***************************************
